library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package reciprocal_pkg is

    --STATE MACHINE
    constant IDLE                       : std_logic_vector(2 downto 0) := "000";
    constant WAIT_FIRST_FULL_12RGB      : std_logic_vector(2 downto 0) := "001";
    constant WAIT_FIRST_FULL_12MASK     : std_logic_vector(2 downto 0) := "010";
    constant WAIT_DONE_PROCESS_1ROWMASK : std_logic_vector(2 downto 0) := "011";
    constant WAIT_DONE_CHANGE_1ROWRGB   : std_logic_vector(2 downto 0) := "100";
    constant WAIT_DONE_SENDING_1_FIFO   : std_logic_vector(2 downto 0) := "101";
    constant RECHARGE_n_NEW_PROCESS     : std_logic_vector(2 downto 0) := "110";




  
  type lut_type is array (1 to 255) of unsigned(31 downto 0);
  constant recip_table : lut_type := (
    1 => x"00010000",
    2 => x"00008000",
    3 => x"00005555",
    4 => x"00004000",
    5 => x"00003333",
    6 => x"00002AAB",
    7 => x"00002492",
    8 => x"00002000",
    9 => x"00001C72",
   10 => x"0000199A",
   11 => x"00001746",
   12 => x"00001555",
   13 => x"000013B1",
   14 => x"00001249",
   15 => x"00001111",
   16 => x"00001000",
   17 => x"00000F0F",
   18 => x"00000E39",
   19 => x"00000D79",
   20 => x"00000CCD",
   21 => x"00000C31",
   22 => x"00000BA3",
   23 => x"00000B21",
   24 => x"00000AAB",
   25 => x"00000A3D",
   26 => x"000009D9",
   27 => x"0000097B",
   28 => x"00000925",
   29 => x"000008D4",
   30 => x"00000889",
   31 => x"00000842",
   32 => x"00000800",
   33 => x"000007C2",
   34 => x"00000788",
   35 => x"00000750",
   36 => x"0000071C",
   37 => x"000006EB",
   38 => x"000006BD",
   39 => x"00000690",
   40 => x"00000666",
   41 => x"0000063E",
   42 => x"00000618",
   43 => x"000005F4",
   44 => x"000005D1",
   45 => x"000005B0",
   46 => x"00000591",
   47 => x"00000572",
   48 => x"00000555",
   49 => x"00000539",
   50 => x"0000051F",
   51 => x"00000505",
   52 => x"000004EC",
   53 => x"000004D5",
   54 => x"000004BE",
   55 => x"000004A8",
   56 => x"00000492",
   57 => x"0000047E",
   58 => x"0000046A",
   59 => x"00000457",
   60 => x"00000444",
   61 => x"00000432",
   62 => x"00000421",
   63 => x"00000410",
   64 => x"00000400",
   65 => x"000003F0",
   66 => x"000003E1",
   67 => x"000003D2",
   68 => x"000003C4",
   69 => x"000003B6",
   70 => x"000003A8",
   71 => x"0000039B",
   72 => x"0000038E",
   73 => x"00000382",
   74 => x"00000376",
   75 => x"0000036A",
   76 => x"0000035E",
   77 => x"00000353",
   78 => x"00000348",
   79 => x"0000033E",
   80 => x"00000333",
   81 => x"00000329",
   82 => x"0000031F",
   83 => x"00000316",
   84 => x"0000030C",
   85 => x"00000303",
   86 => x"000002FA",
   87 => x"000002F1",
   88 => x"000002E9",
   89 => x"000002E0",
   90 => x"000002D8",
   91 => x"000002D0",
   92 => x"000002C8",
   93 => x"000002C1",
   94 => x"000002B9",
   95 => x"000002B2",
   96 => x"000002AB",
   97 => x"000002A4",
   98 => x"0000029D",
   99 => x"00000296",
  100 => x"0000028F",
  101 => x"00000289",
  102 => x"00000283",
  103 => x"0000027C",
  104 => x"00000276",
  105 => x"00000270",
  106 => x"0000026A",
  107 => x"00000264",
  108 => x"0000025F",
  109 => x"00000259",
  110 => x"00000254",
  111 => x"0000024E",
  112 => x"00000249",
  113 => x"00000244",
  114 => x"0000023F",
  115 => x"0000023A",
  116 => x"00000235",
  117 => x"00000230",
  118 => x"0000022B",
  119 => x"00000227",
  120 => x"00000222",
  121 => x"0000021E",
  122 => x"00000219",
  123 => x"00000215",
  124 => x"00000211",
  125 => x"0000020C",
  126 => x"00000208",
  127 => x"00000204",
  128 => x"00000200",
  129 => x"000001FC",
  130 => x"000001F8",
  131 => x"000001F4",
  132 => x"000001F0",
  133 => x"000001ED",
  134 => x"000001E9",
  135 => x"000001E5",
  136 => x"000001E2",
  137 => x"000001DE",
  138 => x"000001DB",
  139 => x"000001D7",
  140 => x"000001D4",
  141 => x"000001D1",
  142 => x"000001CE",
  143 => x"000001CA",
  144 => x"000001C7",
  145 => x"000001C4",
  146 => x"000001C1",
  147 => x"000001BE",
  148 => x"000001BB",
  149 => x"000001B8",
  150 => x"000001B5",
  151 => x"000001B2",
  152 => x"000001AF",
  153 => x"000001AC",
  154 => x"000001AA",
  155 => x"000001A7",
  156 => x"000001A4",
  157 => x"000001A1",
  158 => x"0000019F",
  159 => x"0000019C",
  160 => x"0000019A",
  161 => x"00000197",
  162 => x"00000195",
  163 => x"00000192",
  164 => x"00000190",
  165 => x"0000018D",
  166 => x"0000018B",
  167 => x"00000188",
  168 => x"00000186",
  169 => x"00000184",
  170 => x"00000182",
  171 => x"0000017F",
  172 => x"0000017D",
  173 => x"0000017B",
  174 => x"00000179",
  175 => x"00000176",
  176 => x"00000174",
  177 => x"00000172",
  178 => x"00000170",
  179 => x"0000016E",
  180 => x"0000016C",
  181 => x"0000016A",
  182 => x"00000168",
  183 => x"00000166",
  184 => x"00000164",
  185 => x"00000162",
  186 => x"00000160",
  187 => x"0000015E",
  188 => x"0000015D",
  189 => x"0000015B",
  190 => x"00000159",
  191 => x"00000157",
  192 => x"00000155",
  193 => x"00000154",
  194 => x"00000152",
  195 => x"00000150",
  196 => x"0000014E",
  197 => x"0000014D",
  198 => x"0000014B",
  199 => x"00000149",
  200 => x"00000148",
  201 => x"00000146",
  202 => x"00000144",
  203 => x"00000143",
  204 => x"00000141",
  205 => x"00000140",
  206 => x"0000013E",
  207 => x"0000013D",
  208 => x"0000013B",
  209 => x"0000013A",
  210 => x"00000138",
  211 => x"00000137",
  212 => x"00000135",
  213 => x"00000134",
  214 => x"00000132",
  215 => x"00000131",
  216 => x"0000012F",
  217 => x"0000012E",
  218 => x"0000012D",
  219 => x"0000012B",
  220 => x"0000012A",
  221 => x"00000129",
  222 => x"00000127",
  223 => x"00000126",
  224 => x"00000125",
  225 => x"00000123",
  226 => x"00000122",
  227 => x"00000121",
  228 => x"0000011F",
  229 => x"0000011E",
  230 => x"0000011D",
  231 => x"0000011C",
  232 => x"0000011A",
  233 => x"00000119",
  234 => x"00000118",
  235 => x"00000117",
  236 => x"00000116",
  237 => x"00000115",
  238 => x"00000113",
  239 => x"00000112",
  240 => x"00000111",
  241 => x"00000110",
  242 => x"0000010F",
  243 => x"0000010E",
  244 => x"0000010D",
  245 => x"0000010B",
  246 => x"0000010A",
  247 => x"00000109",
  248 => x"00000108",
  249 => x"00000107",
  250 => x"00000106",
  251 => x"00000105",
  252 => x"00000104",
  253 => x"00000103",
  254 => x"00000102",
  255 => x"00000101"
  );

end package reciprocal_pkg;